module pixels

pub struct Vector2 {
pub:
	x int
	y int
}